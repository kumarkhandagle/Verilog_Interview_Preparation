module top(input a,b,c,d, input [1:0] sel, output reg y);
  
//////////////////Start Writing your code from here ///////////  

  
  
  
  
  
  
  
  
  
  
  
  
///////////////////End your code above this line /////////////  
endmodule