module top(input clk, input rst, output reg r,y,g);

////////////Start Writing your code here///////////////

  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
 /////////////////////End your code here //////////////////// 
endmodule