module uart_clk (
input clk,    ///Board Clock Pin
input start,   //// Start providing clock to UART Module
output reg clkout  //// Desired clock  source for UART Module
);
  
////////////Start Writing your code here /////////////////

  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
 
///////////////////Finish your code here//////////////////////////  
endmodule