`timescale 1ns / 1ps

module top(
input wen, /// Write Enable
input clk,
  input [6:0] addr, /// Address
  input [7:0] din,	/// Data in
  output reg [7:0] dout  /// Data out
);
  
////////////////Start Writing your code here //////////  


  
  
  
  
  
  
  
  
  
  
  
///////////////////Finish your code here ///////////////  
endmodule