module top(
input clk, 			///Input Clock Source 10 nSec
output reg clkout); ////Clkout declare as temp
  
integer temp;  ///////Counter Variable for Clock Generation
  
initial begin   ////Initialization of temp, clkout
  	temp = 0;
    clkout = 0;
end
  
//////Start writing your Logic from here  

  
  
  
  
  
/////End Your Code Here  
endmodule